module PC(Clock , PCin, PCout);
    input [31:0] PCin;
    input Clock;
    output reg [31:0] PCout;

endmodule
