module PC();
    


endmodule